`timescale 1ns/1ps

module tb_asm():
    

endmodule