module PPU_asm()


endmodule