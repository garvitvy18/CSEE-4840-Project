module PPU()


endmodule